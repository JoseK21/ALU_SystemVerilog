module Shift_circular_right #(parameter N = 3)(input logic [N-1:0] a, b, output logic [N-1:0] d8);
	reg signed [N-1:0] temp;
	assign temp = a;
	
	
endmodule
